library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

entity nexys3_sseg_driver is
    port( 
		MY_CLK 	: in  STD_LOGIC;
		DIGIT0  : in  STD_LOGIC_VECTOR (7 downto 0);
		DIGIT1  : in  STD_LOGIC_VECTOR (7 downto 0);
		DIGIT2  : in  STD_LOGIC_VECTOR (7 downto 0);
		DIGIT3  : in  STD_LOGIC_VECTOR (7 downto 0);
		SSEG_CA : out STD_LOGIC_VECTOR (7 downto 0);
		SSEG_AN : out STD_LOGIC_VECTOR (3 downto 0)
	);
end nexys3_sseg_driver;

architecture Behavioral of nexys3_sseg_driver is

	signal refrclk	: STD_LOGIC := '0';
	signal ch_sel	: integer range 0 to 3 := 0;
	signal counter	: integer range 0 to 124999 := 0;

begin

FREQ_DIV: process (MY_CLK) begin
	if rising_edge(MY_CLK) then
		if (counter = 124999) then -- 400Hz Clock, each SSEG will be refreshed with a freq 100Hz 
			refrclk <= not refrclk;
			counter <= 0;
		else
			counter <= counter + 1;
		end if;
	end if;
end process;
    
process(refrclk) begin
	if rising_edge(refrclk) then
		if (ch_sel = 3) then
			ch_sel <= 0;
		else
			ch_sel <= ch_sel + 1;
		end if;
	end if;
end process;
	
with ch_sel select
	SSEG_AN <= 
		"0111" when 0,
		"1011" when 1,
		"1101" when 2,
		"1110" when 3;

with ch_sel select
	SSEG_CA <= 
		DIGIT0 when 0,
		DIGIT1 when 1,
		DIGIT2 when 2,
		DIGIT3 when 3;

end Behavioral;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;


entity vgadriver is
    Port ( 		
	            seviye : in integer;
					a1 : in integer;
					a2 : in integer;
					b1 : in integer;
					b2 : in integer;
					
					x11:in integer;
					x12:in integer;
					y11:in integer;
					y12:in integer;
					
					
					x21:in integer;
					x22:in integer;
					y21:in integer;
					y22:in integer;
					
					
					x31:in integer;
					x32:in integer;
					y31:in integer;
					y32:in integer;
					
					x41:in integer;
					x42:in integer;
					y41:in integer;
					y42:in integer;
					
					x51:in integer;
					x52:in integer;
					y51:in integer;
					y52:in integer;
					
					x61:in integer;
					x62:in integer;
					y61:in integer;
					y62:in integer;
					
					x71:in integer;
					x72:in integer;
					y71:in integer;
					y72:in integer;
              
               x81:in integer;
					x82:in integer;
					y81:in integer;
					y82:in integer;
					
					
              clk : in  STD_LOGIC;
				  nreset : in std_logic;
              hsync : out  STD_LOGIC;
              vsync : out  STD_LOGIC;
              RGB : out std_logic_vector(7 downto 0)
            );
end vgadriver;

architecture Behavioral of vgadriver is
    signal renktutucu : integer :=0;
    signal vcount : integer := 0;
    signal temp : STD_LOGIC := '0';
	 signal t: std_logic;
	 signal counterresult : std_logic_vector(7 downto 0) :="00000000";
	 signal counter1 : integer range  0 to 1 :=0;
	 signal hcount : integer := 0;
	 signal screenlast : std_logic :='1';
	 
	 
	 
	 type won is array (0 to 55) of std_logic_vector(0 to 279);
  constant screenwon: won:=(("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111",
"1111100000111111111111111111100000111111111111111111000000000000111111111111111111111100001111111111111111111110000011111111111111111111111000001111111111111111111000001111111111111111111100000111111111000011111111111110000011111111111111111111000011111111111111110000011111111111",
"1111100000011111111111111111100000111111111111111000000000000000000111111111111111111000001111111111111111111110000011111111111111111111111000001111111111111111111000000111111111111111111100000111111110000011111111111100000000111111111111111111000001111111111111110000011111111111",
"1111100000011111111111111111000000111111111111100000000000000000000001111111111111111000001111111111111111111110000011111111111111111111111000000111111111111111110000000111111111111111111000000111111110000011111111111100000000111111111111111111000001111111111111110000011111111111",
"1111110000001111111111111111000000111111111111000000000000000000000000111111111111111000001111111111111111111110000011111111111111111111111000000111111111111111110000000111111111111111111000000111111110000011111111111100000000011111111111111111000001111111111111110000011111111111",
"1111110000001111111111111110000001111111111110000000000011110000000000011111111111111000001111111111111111111110000011111111111111111111111000000111111111111111110000000011111111111111111000000111111110000011111111111100000000001111111111111111000001111111111111110000011111111111",
"1111111000000111111111111110000001111111111100000000111111111110000000001111111111111000001111111111111111111110000011111111111111111111111100000111111111111111110000000011111111111111111000001111111110000011111111111100000000001111111111111111000001111111111111110000011111111111",
"1111111000000111111111111100000011111111111000000011111111111111100000000111111111111000001111111111111111111110000011111111111111111111111100000011111111111111100000000011111111111111110000001111111110000011111111111100000000000111111111111111000001111111111111110000011111111111",
"1111111100000011111111111100000011111111110000000111111111111111110000000111111111111000001111111111111111111110000011111111111111111111111100000011111111111111100000000001111111111111110000001111111110000011111111111100000000000111111111111111000001111111111111110000011111111111",
"1111111100000011111111111000000111111111110000001111111111111111111000000011111111111000001111111111111111111110000011111111111111111111111110000011111111111111100000000001111111111111110000011111111110000011111111111100000100000011111111111111000001111111111111110000011111111111",
"1111111110000001111111111000000111111111100000011111111111111111111100000011111111111000001111111111111111111110000011111111111111111111111110000001111111111111100000000001111111111111110000011111111110000011111111111100000100000011111111111111000001111111111111110000011111111111",
"1111111110000001111111110000001111111111100000011111111111111111111100000001111111111000001111111111111111111110000011111111111111111111111110000001111111111111000001000001111111111111100000011111111110000011111111111100000110000001111111111111000001111111111111110000011111111111",
"1111111111000000111111110000001111111111000000111111111111111111111110000001111111111000001111111111111111111110000011111111111111111111111110000001111111111111000001000000111111111111100000111111111110000011111111111100000110000001111111111111000001111111111111110000011111111111",
"1111111111000000111111100000011111111111000000111111111111111111111110000001111111111000001111111111111111111110000011111111111111111111111111000001111111111111000001000000111111111111100000111111111110000011111111111100000111000000111111111111000001111111111111110000011111111111",
"1111111111100000111111100000011111111111000000111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111000000111111111111000011100000111111111111100000111111111110000011111111111100000111000000011111111111000001111111111111110000011111111111",
"1111111111100000011111000000111111111111000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111000000111111111110000011100000111111111111000000111111111110000011111111111100000111100000011111111111000001111111111111110000011111111111",
"1111111111110000011111000000111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111100000111111111110000011100000011111111111000001111111111110000011111111111100000111100000001111111111000001111111111111110000011111111111",
"1111111111110000001110000001111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111100000111111111110000011110000011111111111000001111111111110000011111111111100000111110000001111111111000001111111111111110000011111111111",
"1111111111111000001110000001111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111100000011111111110000111110000011111111110000001111111111110000011111111111100000111111000000111111111000001111111111111110000011111111111",
"1111111111111000000110000011111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111100000011111111100000111110000001111111110000011111111111110000011111111111100000111111000000111111111000001111111111111110000011111111111",
"1111111111111100000100000011111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111110000011111111100000111110000001111111110000011111111111110000011111111111100000111111100000011111111000001111111111111110000011111111111",
"1111111111111100000000000111111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111110000001111111100000111111000001111111110000011111111111110000011111111111100000111111100000011111111000001111111111111110000011111111111",
"1111111111111110000000000111111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111110000001111111100001111111000001111111100000011111111111110000011111111111100000111111110000001111111000001111111111111110000011111111111",
"1111111111111110000000001111111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111111000001111111000001111111000000111111100000111111111111110000011111111111100000111111110000001111111000001111111111111110000011111111111",
"1111111111111111000000001111111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111111000001111111000001111111100000111111100000111111111111110000011111111111100000111111111000000111111000001111111111111110000011111111111",
"1111111111111111000000011111111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111111000000111111000001111111100000111111100000111111111111110000011111111111100000111111111000000011111000001111111111111110000011111111111",
"1111111111111111100000011111111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111111000000111111000011111111100000011111000001111111111111110000011111111111100000111111111100000011111000001111111111111110000011111111111",
"1111111111111111100000111111111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111111100000111110000011111111100000011111000001111111111111110000011111111111100000111111111110000001111000001111111111111110000011111111111",
"1111111111111111100000111111111111111110000001111111111111111111111111000000111111111000001111111111111111111110000011111111111111111111111111111100000111110000011111111110000011111000001111111111111110000011111111111100000111111111110000001111000001111111111111110000011111111111",
"1111111111111111100000111111111111111110000001111111111111111111111110000001111111111000000111111111111111111110000011111111111111111111111111111100000011110000011111111110000011111000001111111111111110000011111111111100000111111111111000000111000001111111111111110000011111111111",
"1111111111111111100000111111111111111111000000111111111111111111111110000001111111111000000111111111111111111110000011111111111111111111111111111110000011110000111111111110000001110000011111111111111110000011111111111100000111111111111000000111000001111111111111110000011111111111",
"1111111111111111100000111111111111111111000000111111111111111111111110000001111111111000000111111111111111111100000011111111111111111111111111111110000011100000111111111110000001110000011111111111111110000011111111111100000111111111111100000011000001111111111111111000011111111111",
"1111111111111111100000111111111111111111000000111111111111111111111100000011111111111000000111111111111111111100000011111111111111111111111111111110000011100000111111111111000001110000011111111111111110000011111111111100000111111111111100000011000001111111111111111111111111111111",
"1111111111111111100000111111111111111111100000011111111111111111111100000011111111111100000011111111111111111100000111111111111111111111111111111110000001100000111111111111000001110000111111111111111110000011111111111100000111111111111110000001000001111111111111111111111111111111",
"1111111111111111100000111111111111111111100000001111111111111111111000000011111111111100000011111111111111111000000111111111111111111111111111111111000001100001111111111111000000100000111111111111111110000011111111111100000111111111111110000001000001111111111111111111111111111111",
"1111111111111111100000111111111111111111110000001111111111111111110000000111111111111100000001111111111111111000000111111111111111111111111111111111000001000001111111111111100000100000111111111111111110000011111111111100000111111111111111000000000001111111111111111111111111111111",
"1111111111111111100000111111111111111111110000000011111111111111100000001111111111111110000000111111111111110000001111111111111111111111111111111111000000000001111111111111100000100000111111111111111110000011111111111100000111111111111111000000000001111111111111110000011111111111",
"1111111111111111100000111111111111111111111000000001111111111111000000001111111111111110000000011111111111000000001111111111111111111111111111111111100000000001111111111111100000000001111111111111111110000011111111111100000111111111111111100000000001111111111111100000001111111111",
"1111111111111111100000111111111111111111111100000000001111111000000000011111111111111111000000000011111100000000011111111111111111111111111111111111100000000011111111111111100000000001111111111111111110000011111111111100000111111111111111110000000001111111111111100000001111111111",
"1111111111111111100000111111111111111111111110000000000000000000000000111111111111111111100000000000000000000000111111111111111111111111111111111111100000000011111111111111110000000001111111111111111110000011111111111100000111111111111111110000000001111111111111100000001111111111",
"1111111111111111100000111111111111111111111111000000000000000000000011111111111111111111110000000000000000000001111111111111111111111111111111111111100000000011111111111111110000000011111111111111111110000011111111111100000111111111111111111000000001111111111111100000001111111111",
"1111111111111111100000111111111111111111111111110000000000000000000111111111111111111111111100000000000000000111111111111111111111111111111111111111110000000011111111111111110000000011111111111111111110000011111111111100000111111111111111111000000001111111111111100000001111111111",
"1111111111111111100000111111111111111111111111111100000000000000111111111111111111111111111111000000000000011111111111111111111111111111111111111111110000000111111111111111111000000011111111111111111110000011111111111100000111111111111111111110000011111111111111110000011111111111",
"1111111111111111111111111111111111111111111111111111111000001111111111111111111111111111111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"));

	 
	 
	 
	 begin

    freqprocess : process(clk,nreset)
    begin
	 if(nreset ='1') then
	 temp <= '0';
        elsif(rising_edge(clk)) then
            if(counter1 = 1) then
				temp <= not temp;
				counter1 <=0;
				else
				counter1 <= counter1 + 1;
				end if;
				end if;
				end process;
				t <= temp;
				
				counter : process(t,nreset)
				begin
				 if(nreset ='1') then
				 counterresult <="00000000";
				elsif(rising_edge(t)) then
				
				
				if(counterresult ="11111111" or hcount >=640) then
				counterresult <= "00000000";
				elsif(seviye=1)then
				counterresult <=  "01110011";
				elsif(seviye=2)then
				counterresult <=  "10101010";
				elsif(seviye=3)then
				counterresult <=  "00000000";
				elsif(seviye=4)then
				counterresult <=  "01010011";
				elsif(seviye=5)then
				counterresult <=  "00000000";
				else 
				counterresult <=  "01010101";
				
				end if ;
				
				if(x11<=hcount and hcount<=x12 and vcount<=y12 and y11<=vcount)then
					if(seviye=1) then
					counterresult <= "00111000";
					end if;
					
					if(seviye=2) then
					counterresult <= "00000011";
					end if;
					
					if(seviye=3) then
					counterresult <= "00010110";
					end if;
					
					if(seviye=4) then
					counterresult <= "00000000";
					end if;
					
				
				end if;
				
				if(x21<=hcount and hcount<=x22 and y21<= vcount and vcount<=y22)then
				
					if(seviye=1) then
					counterresult <= "00111000";
					end if;
					
					if(seviye=2) then
					counterresult <= "00000011";
					end if;
					
					if(seviye=3) then
					counterresult <= "00010110";
					end if;
					
					if(seviye=4) then
					counterresult <= "00000000";
					end if;
				
				end if;
				
				if(x31<=hcount and hcount<=x32 and y31<=vcount and vcount<=y32)then
				
				
					if(seviye=1) then
					counterresult <= "00111000";
					end if;
					
					if(seviye=2) then
					counterresult <= "00000011";
					end if;
					
					if(seviye=3) then
					counterresult <= "00010110";
					end if;
					
					if(seviye=4) then
					counterresult <= "00000000";
					end if;
				
				
				end if;
				
				if(x41<=hcount and hcount<=x42 and y41<=vcount and vcount<=y42)then
				
				
					if(seviye=1) then
					counterresult <= "00111000";
					end if;
					
					if(seviye=2) then
					counterresult <= "00000011";
					end if;
					
					if(seviye=3) then
					counterresult <= "00010110";
					end if;
					
					if(seviye=4) then
					counterresult <= "00000000";
					end if;
				
				
				end if;
				
				if(x51<=hcount and hcount<=x52 and vcount>=y51 and vcount<=y52)then
				
				
					if(seviye=1) then
					counterresult <= "00111000";
					end if;
					
					if(seviye=2) then
					counterresult <= "00000011";
					end if;
					
					if(seviye=3) then
					counterresult <= "00010110";
					end if;
					
					if(seviye=4) then
					counterresult <= "00000000";
					end if;
					
					
				end if;
				
				if(x61<=hcount and hcount<=x62 and y61<=vcount and vcount<=y62)then
				
					if(seviye=1) then
					counterresult <= "00111000";
					end if;
					
					if(seviye=2) then
					counterresult <= "00000011";
					end if;
					
					if(seviye=3) then
					counterresult <= "00010110";
					end if;
					
					if(seviye=4) then
					counterresult <= "00000000";
					end if;
				
				
				end if;
				
				if(x71<=hcount and hcount<=x72 and vcount<=y72 and y71<=vcount) then
				
				
					if(seviye=1) then
					counterresult <= "00111000";
					end if;
					
					if(seviye=2) then
					counterresult <= "00000011";
					end if;
					
					if(seviye=3) then
					counterresult <= "00010110";
					end if;
					
					if(seviye=4) then
					counterresult <= "00000000";
					end if;
				
				
				end if;
--Burda belli aralklarda kutucuk yaptm.
-- odul kutusunu belirledim
				if(x81<=hcount and hcount<=x82 and vcount<=y82 and y81<=vcount) then
				counterresult <= "11111000";
				end if;
				
				
				if(a1<=hcount and hcount<=a2 and b1<=vcount and vcount<=b2 and seviye<5)then
				counterresult <= "11000000";
				
				end if;
				if(seviye=5) then
				
--				if(vcount<240 or vcount>247 or hcount<300 or hcount>344) then
--				counterresult <= "00000000";
--				elsif(screenwon(vcount-240)(hcount-300)='0') then
--				counterresult <= "11100000";
--				else
--				counterresult <= "00000000";
--				end if;
--				
				if (vcount>=212 and vcount<=267 and hcount>=180 and hcount<=459)then
					if(screenwon(vcount-212)(hcount-180)='0') then
						counterresult <= "00000011";
					else
						counterresult <= "11111111";
					end if;
					else 
					 counterresult <= "11111111";
				end if;
				end if;				
				
				
				
				end if;
				end process;
				
				
				
				gulkah : process(t,nreset)
				begin
				 if(nreset ='1') then
				 hcount <= 0;
				 vcount <= 0;
            elsif(t = '1' and t' event) then         -- Happens at 25MHz (50MHz / 2)

                -- Reset the counter if column/line finished or increment it
                if(hcount = 799) then
                    hcount <= 0;
                    if vcount = 521 then
                        vcount <= 0;
                    else
                        vcount <= vcount + 1;
                    end if;
                else
                    hcount <= hcount + 1;
                end if;
               end if;
					end process;
					
					
                -- Send a pulse of vsync to start a new column
					 
                kah : process(t,nreset)
					 begin
					  if(nreset ='1') then
					  vsync <= '0';
					  hsync <= '0';
					 elsif(rising_edge(t)) then
					 if vcount >= 490 and vcount < 492 then
                    vsync <= '0';
                else
                    vsync <= '1';	
                end if;

                -- Send a pulse of hsync to start a new line
                if hcount >= 656 and hcount < 752 then
                    hsync <= '0';
                else
                    hsync <= '1';
                end if;
                  end if;
						end process;
                -- If pixel time, draw something
					 
					 
					 
					 
                disp : process(t,nreset)
					 begin
					  if(nreset ='1') then
					  RGB <= "00000000";
					 elsif(rising_edge(t)) then
					 if (hcount < 640 and vcount < 480)  then
                   
						 RGB <= counterresult;
                else
                   RGB <="00000000";
                end if;
					 end if;
					 end process;
           

end Behavioral;
LIBRARY ieee ;
 USE ieee.std_logic_1164.all ;
 
 USE ieee.std_logic_arith.all ;
 USE ieee.std_logic_unsigned.all;
 
 --buradansonra 
 


entity seviye_to_seven_segment is
port(d: in integer; s: out std_logic_vector(6 downto 0));
end seviye_to_seven_segment;

architecture dataflow of seviye_to_seven_segment is 

begin 

s <="1000000" when d=1 else
"1111001" when d=2 else 
"0100100" when d=3 else 
"0110000" when d=4 else
"0011001" when d=5 else 
"0010010" when d=6 else 
"0000010" when d=7 else 
"1111000" when d=8 else 
"0000000" when d=9 else 
"0010000" when d=10 else 
"1111111"; 

end dataflow; 

LIBRARY ieee ;
 USE ieee.std_logic_1164.all ;
 
 USE ieee.std_logic_arith.all ;
 USE ieee.std_logic_unsigned.all;
 
 
 --buradan oce
 
 
 
 
 
 entity ee240_vgadriver is
  port (right1 : in std_logic :='0';
  left1 : in std_logic :='0';
  up1 : in std_logic :='0';
  down1 : in std_logic :='0';
  nreset: in std_logic;
  board_clk: in std_logic;
  vsync: out std_logic;
  hsync: out std_logic;
  red: out std_logic_vector(2 downto 0);
  green: out std_logic_vector(2 downto 0);
  blue: out std_logic_vector(1 downto 0);
  CA : out STD_LOGIC_VECTOR (7 downto 0);
  AN : out STD_LOGIC_VECTOR (3 downto 0));
 end ee240_vgadriver;
 architecture arch_vga_driver of ee240_vgadriver is
 component gullukkahraman
  Port ( 	seviye:in integer;
           a1 : in integer;
				a2 : in integer;
				b1 : in integer;
				b2 : in integer;
				
				x11:in integer;
					x12:in integer;
					y11:in integer;
					y12:in integer;
					
					
					x21:in integer;
					x22:in integer;
					y21:in integer;
					y22:in integer;
					
					
					x31:in integer;
					x32:in integer;
					y31:in integer;
					y32:in integer;
					
					x41:in integer;
					x42:in integer;
					y41:in integer;
					y42:in integer;
					
					x51:in integer;
					x52:in integer;
					y51:in integer;
					y52:in integer;
					
					x61:in integer;
					x62:in integer;
					y61:in integer;
					y62:in integer;
					
					x71:in integer;
					x72:in integer;
					y71:in integer;
					y72:in integer;
					
					x81:in integer;
					x82:in integer;
					y81:in integer;
					y82:in integer;
				
				
				
				clk : in  STD_LOGIC;
				nreset : in std_logic;
            hsync : out  STD_LOGIC;
            vsync : out  STD_LOGIC;
            RGB : out std_logic_vector(7 downto 0));
 end component;
  for all : gullukkahraman use entity work.vgadriver(Behavioral);
  
  --buuuu
  component seviyedensevensegmente
  Port (  d : in integer;
				
           s : out std_logic_vector(6 downto 0));
 end component;

  for all : seviyedensevensegmente use entity work.seviye_to_seven_segment(dataflow);
  
  component nexy			
			port( 
		MY_CLK 	: in  STD_LOGIC;
		DIGIT0  : in  STD_LOGIC_VECTOR (7 downto 0);
		DIGIT1  : in  STD_LOGIC_VECTOR (7 downto 0);
		DIGIT2  : in  STD_LOGIC_VECTOR (7 downto 0);
		DIGIT3  : in  STD_LOGIC_VECTOR (7 downto 0);
		SSEG_CA : out STD_LOGIC_VECTOR (7 downto 0);
		SSEG_AN : out STD_LOGIC_VECTOR (3 downto 0)
	);
	end component;
	for all : nexy use entity work.nexys3_sseg_driver (Behavioral);
  
  
  --buuuu
  
  
  
  
  
  signal RGB : std_logic_vector(7 downto 0);
  signal controller : integer range 0 to 4168799:=0 ;
  signal controller2 : integer range 0 to 10000000:=0 ;
  signal turp : integer range 0 to 416799 :=0;
  signal seviye : integer range 1 to 10 :=1; 
  signal a1 : integer range 0 to 640 :=5;
  signal a2 : integer range 0 to 640 :=15;
  signal b1 : integer range 0 to 480 :=235;
  signal b2 : integer range 0 to 480 :=250;
  
  signal x11 : integer range 0 to 639 :=170;
  signal x12 : integer range 0 to 639 :=180;
  signal y11 : integer range 0 to 479 :=0;
  signal y12 : integer range 0 to 479 :=120;
  
  signal x21 : integer range 0 to 639 :=240;
  signal x22 : integer range 0 to 639 :=250;
  signal y21 : integer range 0 to 479 :=339;
  signal y22 : integer range 0 to 479 :=479;
  
  signal x31 : integer range 0 to 639 :=290;
  signal x32 : integer range 0 to 639 :=300;
  signal y31 : integer range 0 to 479 :=150;
  signal y32 : integer range 0 to 479 :=280;
  
  signal x41 : integer range 0 to 639 :=360;
  signal x42 : integer range 0 to 639 :=370;
  signal y41 : integer range 0 to 479 :=0;
  signal y42 : integer range 0 to 479 :=100;
  
  signal x51 : integer range 0 to 639 :=440;
  signal x52 : integer range 0 to 639 :=450;
  signal y51 : integer range 0 to 479 :=280;
  signal y52 : integer range 0 to 479 :=479;
  
  signal x61 : integer range 0 to 639 :=500;
  signal x62 : integer range 0 to 639 :=510;
  signal y61 : integer range 0 to 479 :=0;
  signal y62 : integer range 0 to 479 :=170;
  
  signal x71 : integer range 0 to 639 :=540;
  signal x72 : integer range 0 to 639 :=550;
  signal y71 : integer range 0 to 479 :=200;
  signal y72 : integer range 0 to 479 :=330;
  
  -- yakalamak istedi sey 
  signal x81 : integer range 0 to 639 :=560;
  signal x82 : integer range 0 to 639 :=565;
  signal y81 : integer range 0 to 479 :=110;
  signal y82 : integer range 0 to 479 :=115;
 
  signal tempa1 : integer range 0 to 640 :=5;
  signal tempa2 : integer range 0 to 640 :=15;
  signal tempb1 : integer range 0 to 480 :=235;
  signal tempb2 : integer range 0 to 480 :=250;
  
 
 
  signal c : integer range 0 to 640 ;
  signal d : integer range 0 to 640 ;
  signal kaykon1 : integer range 0 to 1 :=0;
  signal kaykon2 : std_logic :='0';
  signal kaykon3 : std_logic :='1';
  signal kaykon4 : std_logic :='1';
  signal kaykon5 : std_logic :='0';
  signal kaykon6 : std_logic :='1';
  signal kaykon7 : std_logic :='0';
  
  
  signal tempy11 : integer range 0 to 479 :=0;
  signal tempy12 : integer range 0 to 479 :=120;
  signal tempy21 : integer range 0 to 479 :=339;
  signal tempy22 : integer range 0 to 479 :=479;
  signal tempy31 : integer range 0 to 479 :=150;
  signal tempy32 : integer range 0 to 479 :=280;
  signal tempy41 : integer range 0 to 479 :=0;
  signal tempy42 : integer range 0 to 479 :=100;
  signal tempy51 : integer range 0 to 479 :=280;
  signal tempy52 : integer range 0 to 479 :=479;
  signal tempy61 : integer range 0 to 479 :=0;
  signal tempy62 : integer range 0 to 479 :=170;
  signal tempy71 : integer range 0 to 479 :=200;
  signal tempy72 : integer range 0 to 479 :=330;
  signal tempx81 : integer range 0 to 639 :=0;
  signal tempx82 : integer range 0 to 639 :=0;
  signal tempy81 : integer range 0 to 639 :=0;
  signal tempy82 : integer range 0 to 639 :=0;
  signal ss : std_logic_vector(6 downto 0);
  signal minnos : std_logic_vector(7 downto 0);
  signal hatasayisi : integer range 0 to 10 :=1;
  signal kk : std_logic_vector(6 downto 0);
  signal minnos2 : std_logic_vector(7 downto 0);
  signal temphatasayisi : integer range 0 to 10 :=1;
  

  
 begin
 		
					 caz5 : process(board_clk)
						begin
						
						
						if(board_clk' event and board_clk='1') then
						
						
						
						if(right1='1' and a1<629) then
						
						tempa1<=a1+1;
						tempa2<=a2+1;
						
						
						end if;
						
						
						if(left1='1' and a1>0) then
						
						tempa1<=a1-1;
						tempa2<=a2-1;
						
						
						end if;
						
						if(up1='1' and b1>0) then
						
						tempb1<=b1-1;
						tempb2<=b2-1;
						
						
						end if;
						
						if(down1='1' and b1<469) then
						
						tempb1<=b1+1;
						tempb2<=b2+1;
						
						
						end if;
						
						
						
						------
						
						
														
						
						if(controller<416799)then
						controller <= controller+1;
						end if; 
						if(controller=416799) then
						controller<=0;
						a1<=tempa1;
						b1<=tempb1;
						a2<=tempa2;
						b2<=tempb2;

						x81<=tempx81;
						x82<=tempx82;
						y81<=tempy81;
						y82<=tempy82;

						end if;
						
						
						
						
					 if(controller=0) then
					 tempa1<=a1;
					 tempa2<=a2;									--Her baslangicta temp degerlerini tekrardan a1lere atadim
					 tempb1<=b1;
					 tempb2<=b2;
					 
					  tempx81<=x81;
					  tempx82<=x82;
					  tempy81<=y81;
					  tempy82<=y82;
					  end if;
							
						
						
					  if((a1+10<x11) or (b1>y12) or (a1>x12) or (b1+10<y11))then
					  else
					  temphatasayisi<=hatasayisi+1;
					  tempa1<=5;
					  tempa2<=15;
					  tempb1<=235;
					  tempb2<=250;
					  end if;
					  
					  if((a1+10<x21) or (b1>y22) or (a1>x22) or (b1+10<y21))then
					  else
					  temphatasayisi<=hatasayisi+1;
					  tempa1<=5;
					  tempa2<=15;
					  tempb1<=235;
					  tempb2<=250;
					  end if;
					  
					  
					  if((a1+10<x31) or (b1>y32) or (a1>x32) or (b1+10<y31))then
					  else
					  temphatasayisi<=hatasayisi+1;
					  tempa1<=5;
					  tempa2<=15;
					  tempb1<=235;
					  tempb2<=250;
					  end if;
					  
					  
					  if((a1+10<x41) or (b1>y42) or (a1>x42) or (b1+10<y41))then
					  else
					  temphatasayisi<=hatasayisi+1;
					  tempa1<=5;
					  tempa2<=15;
					  tempb1<=235;
					  tempb2<=250;
					  end if;
					  
					  
					  if((a1+10<x51) or (b1>y52) or (a1>x52) or (b1+10<y51))then
					  else
					  temphatasayisi<=hatasayisi+1;
					  tempa1<=5;
					  tempa2<=15;
					  tempb1<=235;
					  tempb2<=250;
					  end if;
					  
					  
					  if((a1+10<x61) or (b1>y62) or (a1>x62) or (b1+10<y61))then
					  else
					  temphatasayisi<=hatasayisi+1;
					  tempa1<=5;
					  tempa2<=15;
					  tempb1<=235;
					  tempb2<=250;
					  end if;
					  
					  if((a1+10<x71) or (b1>y72) or (a1>x72) or (b1+10<y71))then
					  else
					  temphatasayisi<=hatasayisi+1;
					  tempa1<=5;
					  tempa2<=15;
					  tempb1<=235;
					  tempb2<=250;
					  end if;
					  
					  --burasi hata olanb
					  
				  if(hatasayisi=6)  then
					  
				  seviye<=1;
					  temphatasayisi<=1;
					  
					  tempx81<=5;
					  tempx82<=10;
					  tempy81<=5;
					  tempy82<=10;
					  
					  x81<=560;
					  x82<=565;
					  y81<=110;
					  y82<=115;
					  
					  
					  x11<=170;
					  x12<=180;
					  
					  x21<=240;
					  x22<=250;
					  
					  x31<=225;
					  x32<=235;
					  
					  x41<=300;
					  x42<=310;
					  
					  x51<=440;
					  x52<=450;
					  
					  x61<=500;
					  x62<=510;
					  
					  x71<=540;
					  x72<=550;
					  
					  
					  
					  end if;
					  
					  
					  --hatanin bitiidi

 					  if((a1+10<x81) or (b1>y82) or (a1>x82) or (b1+10<y81))then
					  elsif(seviye=1) then
					  tempx81<=5;
					  tempx82<=10;
					  tempy81<=5;
					  tempy82<=10;
					  
					  x81<=5;
					  x82<=10;
					  y81<=5;
					  y82<=10;
					  seviye<=2;
					  
					  x11<=40;
					  x12<=50;
					  
					  x21<=100;
					  x22<=110;
					  
					  x31<=290;
					  x32<=300;
					  
					  x41<=360;
					  x42<=370;
					  
					  x51<=390;
					  x52<=400;
					  
					  x61<=480;
					  x62<=490;
					  
					  x71<=560;
					  x72<=570;
					  
					  
					  					 					  					  					  
					  					
					  
					  end if;

					 if((a1+10<x81) or (b1>y82) or (a1>x82) or (b1+10<y81))then
					  elsif(seviye=2) then
					  tempx81<=625;
					  tempx82<=630;
					  tempy81<=400;
					  tempy82<=405;
					  
					  x81<=625;
					  x82<=630;
					  y81<=400;
					  y82<=405;				  			
					  seviye<=3;
					  
					  x11<=60;
					  x12<=70;
					  
					  x21<=120;
					  x22<=130;
					  
					  x31<=160;
					  x32<=170;
					  
					  x41<=220;
					  x42<=230;
					  
					  x51<=330;
					  x52<=340;
					  
					  x61<=480;
					  x62<=490;
					  
					  x71<=560;
					  x72<=570;
					  
					  
					 
					  end if;
					  
					  if((a1+10<x81) or (b1>y82) or (a1>x82) or (b1+10<y81))then
					  elsif(seviye=3) then
					  tempx81<=50;
					  tempx82<=55;
					  tempy81<=110;
					  tempy82<=115;
					  
					  x81<=50;
					  x82<=55;
					  y81<=110;
					  y82<=115;				  			
					  seviye<=4;
					  x11<=70;
					  x12<=80;
					  
					  x21<=140;
					  x22<=150;
					  
					  x31<=200;
					  x32<=210;
					  
					  x41<=260;
					  x42<=270;
					  
					  x51<=340;
					  x52<=350;
					  
					  x61<=400;
					  x62<=410;
					  
					  x71<=500;
					  x72<=510;
					  
					 
					  end if;
					  
					  if((a1+10<x81) or (b1>y82) or (a1>x82) or (b1+10<y81))then
					  elsif(seviye=4) then
					  tempx81<=0;
					  tempx82<=0;
					  tempy81<=0;
					  tempy82<=0;
					  
					  x81<=0;
					  x82<=0;
					  y81<=0;
					  y82<=0;				  			
					  seviye<=5;
					  
					  x11<=0;
					  x12<=0;
					  
					  x21<=0;
					  x22<=0;
					  
					  x31<=0;
					  x32<=0;
					  
					  x41<=0;
					  x42<=0;
					  
					  x51<=0;
					  x52<=0;
					  
					  x61<=0;
					  x62<=0;
					  
					  x71<=0;
					  x72<=0;
					  
					 
					  
					 
					  end if;
					  
					  
						
						
						end if;
					 end process;
					 --KESISME SARTLARI BITISI
 
 --DUVARLARIN HAREKET KODUNUN BASLANGICI
 
			kaymalar : process(board_clk)
				begin
				if(board_clk' event and board_clk='1') then
 
				
				if(kaykon1=1) then 
				tempy11<=y11+1;
				tempy12<=y12+1;
				else
				tempy11<=y11-1;
				tempy12<=y12-1;
				end if;
				
				if(tempy12=479) then
				kaykon1<=0;
				tempy11<=y11-1;
				tempy12<=y12-1;
				
				end if;
				
				if(tempy11=1) then
				kaykon1<=1;
				tempy11<=y11+1;
				tempy12<=y12+1;
				
				end if;
				
				
				
				
				
				
				if(kaykon2='1') then 
				tempy21<=y21+1;
				tempy22<=y22+1;
				else
				tempy21<=y21-1;
				tempy22<=y22-1;
				end if;
				
				if(y22=479) then
				kaykon2<='0';
				end if;
				
				if(y21=0) then
				kaykon2<='1';
				end if;
				
				
				
				
				
				
				
				
				if(kaykon3='1') then 
				tempy31<=y31+1;
				tempy32<=y32+1;
				else
				tempy31<=y31-1;
				tempy32<=y32-1;
				end if;
				
				if(y32=479) then
				kaykon3<='0';
				end if;
				
				if(y31=0) then
				kaykon3<='1';
				end if;
				
				
				
				
				
				
				
				if(kaykon4='1') then 
				tempy41<=y41+1;
				tempy42<=y42+1;
				else
				tempy41<=y41-1;
				tempy42<=y42-1;
				end if;
				
				if(y42=479) then
				kaykon4<='0';
				end if;
				
				if(y41=0) then
				kaykon4<='1';
				end if;
				
				
				
				
				
				
				
				if(kaykon5='1') then 
				tempy51<=y51+1;
				tempy52<=y52+1;
				else
				tempy51<=y51-1;
				tempy52<=y52-1;
				end if;
				
				if(y52=479) then
				kaykon5<='0';
				end if;
				
				if(y51=0) then
				kaykon5<='1';
				end if;
				
				
				
				
				
				
				if(kaykon6='1') then 
				tempy61<=y61+1;
				tempy62<=y62+1;
				else
				tempy61<=y61-1;
				tempy62<=y62-1;
				end if;
				
				if(y62=479) then
				kaykon6<='0';
				end if;
				
				if(y61=0) then
				kaykon6<='1';
				end if;
				
				
				
				
				
				
				
				if(kaykon7='1') then 
				tempy71<=y71+1;
				tempy72<=y72+1;
				else
				tempy71<=y71-1;
				tempy72<=y72-1;
				end if;
				
				if(y72=479) then
				kaykon7<='0';
				end if;
				
				if(y71=0) then
				kaykon7<='1';
				end if;
				
				
				
				
				
				
				if(turp>=0) then
				turp<=turp+1;
				end if;
				
				
			
				
				
				if(turp=416799) then
				y11<=tempy11;
				y12<=tempy12; 
				y21<=tempy21;
				y22<=tempy22;
				y31<=tempy31;
				y32<=tempy32;
				y41<=tempy41;
				y42<=tempy42;
				y51<=tempy51;
				y52<=tempy52;
				y61<=tempy61;
				y62<=tempy62;
				y71<=tempy71;
				y72<=tempy72;
				turp<=0;
				hatasayisi<=temphatasayisi;
				end if;
				
				
				
				
				
				
				
				end if;
				end process;
 
 
 
 
 
 --DUVARLARIN HAREKET KODUNUN Bitisi
 
 
 
 
 c<=a1+10;
 d<=b1+10;
 
 
 munir1 : seviyedensevensegmente port map(seviye,ss);
 munir2 : seviyedensevensegmente port map(hatasayisi,kk);
 kapi1 : gullukkahraman port map(seviye,a1,c,b1,d,x11,x12,y11,y12,x21,x22,y21,y22,x31,x32,y31,y32,x41,x42,y41,y42,x51,x52,y51,y52,x61,x62,y61,y62,x71,x72,y71,y72,x81,x82,y81,y82,board_clk,nreset,hsync,vsync,RGB);
 red <= RGB(7 downto 5);
 green <= RGB(4 downto 2);
 blue <= RGB(1 downto 0);
 
 minnos(7)<='1';
 minnos(6 downto 0) <= ss(6 downto 0);
 
 minnos2(7)<='1';
 minnos2(6 downto 0) <= kk(6 downto 0);
 
 
 RESULT : nexy PORT MAP	(board_clk,minnos2,"11111111",minnos,"11000000",CA,AN);	

 end arch_vga_driver;